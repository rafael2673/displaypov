library ieee;
use ieee.std_logic_1164.all;

package TypesPackage is
	type matrix_type is array (0 to 7) of std_logic_vector(7 downto 0);
end package TypesPackage;
