library ieee;
use ieee.std_logic_1164.all;

entity pov is
   port (SW: in  std_logic_vector(3 downto 0);
			KEY: in std_logic_vector(2 downto 0);
                       LEDR, LEDG : out std_logic_vector(7 downto 0));
end pov;

architecture logica of pov is

type matrix_type is array(0 to 7, 0 to 7) of std_logic;

constant zero_pattern : matrix_type := (
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '0', '1', '1', '1', '0', '0' ),
    ( '0', '0', '1', '0', '0', '0', '1', '0' ),
    ( '0', '0', '1', '0', '0', '1', '1', '0' ),
    ( '0', '0', '1', '0', '1', '0', '1', '0' ),
    ( '0', '0', '1', '1', '0', '0', '1', '0' ),
    ( '0', '0', '1', '0', '0', '0', '1', '0' ),
    ( '0', '0', '0', '1', '1', '1', '0', '0' )
);

constant one_pattern : matrix_type := (
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '0', '0', '1', '0', '0', '0' ),
    ( '0', '0', '0', '1', '1', '0', '0', '0' ),
    ( '0', '0', '0', '0', '1', '0', '0', '0' ),
    ( '0', '0', '0', '0', '1', '0', '0', '0' ),
    ( '0', '0', '0', '0', '1', '0', '0', '0' ),
    ( '0', '0', '0', '0', '1', '0', '0', '0' ),
    ( '0', '0', '0', '1', '1', '1', '0', '0' )
);

constant two_pattern : matrix_type := (
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '0', '1', '1', '1', '0', '0' ),
    ( '0', '0', '1', '0', '0', '0', '1', '0' ),
    ( '0', '0', '0', '0', '0', '0', '1', '0' ),
    ( '0', '0', '0', '0', '1', '1', '0', '0' ),
    ( '0', '0', '0', '1', '0', '0', '0', '0' ),
    ( '0', '0', '1', '0', '0', '0', '0', '0' ),
    ( '0', '0', '1', '1', '1', '1', '1', '0' )
);

constant three_pattern : matrix_type := (
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '0', '1', '1', '1', '0', '0' ),
    ( '0', '0', '1', '0', '0', '0', '1', '0' ),
    ( '0', '0', '0', '0', '0', '0', '1', '0' ),
    ( '0', '0', '0', '1', '1', '1', '0', '0' ),
    ( '0', '0', '0', '0', '0', '0', '1', '0' ),
    ( '0', '0', '1', '0', '0', '0', '1', '0' ),
    ( '0', '0', '0', '1', '1', '1', '0', '0' )
);

constant four_pattern : matrix_type := (
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '0', '0', '0', '1', '0', '0' ),
    ( '0', '0', '0', '0', '1', '1', '0', '0' ),
    ( '0', '0', '0', '1', '0', '1', '0', '0' ),
    ( '0', '0', '1', '0', '0', '1', '0', '0' ),
    ( '0', '0', '1', '1', '1', '1', '1', '0' ),
    ( '0', '0', '0', '0', '0', '1', '0', '0' ),
    ( '0', '0', '0', '0', '0', '1', '0', '0' )
);

constant five_pattern : matrix_type := (
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '1', '1', '1', '1', '1', '0' ),
    ( '0', '0', '1', '0', '0', '0', '0', '0' ),
    ( '0', '0', '1', '1', '1', '1', '0', '0' ),
    ( '0', '0', '0', '0', '0', '0', '1', '0' ),
    ( '0', '0', '0', '0', '0', '0', '1', '0' ),
    ( '0', '0', '1', '0', '0', '0', '1', '0' ),
    ( '0', '0', '0', '1', '1', '1', '0', '0' )
);

constant six_pattern : matrix_type := (
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '0', '0', '1', '1', '0', '0' ),
    ( '0', '0', '0', '1', '0', '0', '0', '0' ),
    ( '0', '0', '1', '0', '0', '0', '0', '0' ),
    ( '0', '0', '1', '1', '1', '1', '0', '0' ),
    ( '0', '0', '1', '0', '0', '0', '1', '0' ),
    ( '0', '0', '1', '0', '0', '0', '1', '0' ),
    ( '0', '0', '0', '1', '1', '1', '0', '0' )
);

constant seven_pattern : matrix_type := (
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '1', '1', '1', '1', '1', '0' ),
    ( '0', '0', '0', '0', '0', '0', '1', '0' ),
    ( '0', '0', '0', '0', '0', '1', '0', '0' ),
    ( '0', '0', '0', '0', '1', '0', '0', '0' ),
    ( '0', '0', '0', '1', '0', '0', '0', '0' ),
    ( '0', '0', '0', '1', '0', '0', '0', '0' ),
    ( '0', '0', '0', '1', '0', '0', '0', '0' )
);

constant eight_pattern : matrix_type := (
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '0', '1', '1', '1', '0', '0' ),
    ( '0', '0', '1', '0', '0', '0', '1', '0' ),
    ( '0', '0', '1', '0', '0', '0', '1', '0' ),
    ( '0', '0', '0', '1', '1', '1', '0', '0' ),
    ( '0', '0', '1', '0', '0', '0', '1', '0' ),
    ( '0', '0', '1', '0', '0', '0', '1', '0' ),
    ( '0', '0', '0', '1', '1', '1', '0', '0' )
);

constant nine_pattern : matrix_type := (
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '0', '1', '1', '1', '0', '0' ),
    ( '0', '0', '1', '0', '0', '0', '1', '0' ),
    ( '0', '0', '1', '0', '0', '0', '1', '0' ),
    ( '0', '0', '0', '1', '1', '1', '1', '0' ),
    ( '0', '0', '0', '0', '0', '0', '1', '0' ),
    ( '0', '0', '0', '0', '0', '1', '0', '0' ),
    ( '0', '0', '0', '1', '1', '0', '0', '0' )
);

constant ten_pattern : matrix_type := (
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '0', '1', '1', '0', '0', '0' ),
    ( '0', '0', '0', '0', '0', '1', '0', '0' ),
    ( '0', '0', '0', '1', '1', '1', '0', '0' ),
    ( '0', '0', '1', '0', '0', '1', '0', '0' ),
    ( '0', '0', '0', '1', '1', '1', '1', '0' )
);

constant eleven_pattern : matrix_type := (
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '1', '0', '0', '0', '0', '0' ),
    ( '0', '0', '1', '0', '0', '0', '0', '0' ),
    ( '0', '0', '1', '0', '1', '1', '0', '0' ),
    ( '0', '0', '1', '1', '0', '0', '1', '0' ),
    ( '0', '0', '1', '0', '0', '0', '1', '0' ),
    ( '0', '0', '1', '0', '0', '0', '1', '0' ),
    ( '0', '0', '1', '1', '1', '1', '0', '0' )
);

constant twelve_pattern : matrix_type := (
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '0', '1', '1', '1', '0', '0' ),
    ( '0', '0', '1', '0', '0', '0', '0', '0' ),
    ( '0', '0', '1', '0', '0', '0', '0', '0' ),
    ( '0', '0', '1', '0', '0', '0', '1', '0' ),
    ( '0', '0', '0', '1', '1', '1', '0', '0' )
);

constant thirteen_pattern : matrix_type := (
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '0', '0', '0', '0', '1', '0' ),
    ( '0', '0', '0', '0', '0', '0', '1', '0' ),
    ( '0', '0', '0', '1', '1', '0', '1', '0' ),
    ( '0', '0', '1', '0', '0', '1', '1', '0' ),
    ( '0', '0', '1', '0', '0', '0', '1', '0' ),
    ( '0', '0', '1', '0', '0', '0', '1', '0' ),
    ( '0', '0', '0', '1', '1', '1', '1', '0' )
);

constant fourteen_pattern : matrix_type := (
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '0', '1', '1', '1', '0', '0' ),
    ( '0', '0', '1', '0', '0', '0', '1', '0' ),
    ( '0', '0', '1', '1', '1', '1', '0', '0' ),
    ( '0', '0', '1', '0', '0', '0', '0', '0' ),
    ( '0', '0', '0', '1', '1', '1', '0', '0' )
);

constant fiveteen_pattern : matrix_type := (
    ( '0', '0', '0', '0', '0', '0', '0', '0' ),
    ( '0', '0', '0', '0', '0', '1', '0', '0' ),
    ( '0', '0', '0', '0', '1', '0', '1', '0' ),
    ( '0', '0', '0', '0', '1', '0', '0', '0' ),
    ( '0', '0', '0', '1', '1', '1', '0', '0' ),
    ( '0', '0', '0', '0', '1', '0', '0', '0' ),
    ( '0', '0', '0', '0', '1', '0', '0', '0' ),
    ( '0', '0', '0', '0', '1', '0', '0', '0' )
);

 mux_16x1 is
   port (A: in std_logic_vector(15 downto 0);
			S: in std_logic_vector(3 downto 0);
			saida: out std_logic);
end component;

component mux_8x1 is
   port (A, B, C, D, E, F, G, H: in std_logic;
			S: in std_logic_vector(2 downto 0);
			saida: out std_logic);
end component;

signal saida_mux_8: 

begin

LEDR <= pattern(saida_mux_8);

LEDG <= pattern(0)(saida_mux_8) & pattern(1)(saida_mux_8) & pattern(2)(saida_mux_8) & pattern(3)(saida_mux_8) &
        pattern(4)(saida_mux_8) & pattern(5)(saida_mux_8) & zero_pattern(6)(saida_mux_8) & pattern(7)(saida_mux_8);

end logica;